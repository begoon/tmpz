module main

fn main() {
	s := 'abc'
	b := s.clone()
	println('s: ${s}, b: ${b}')
}
