module main

fn main() {
	s := 'abc'
	b := s
	println('s: ${s}, b: ${b}')
}
